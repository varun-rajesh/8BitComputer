module d_ff();

endmodule

module jk_ff();

endmodule
